module vamk

// @TODO: Use a map ?
// Long list of tokens
const token_str_ifeq = 'ifeq'
const token_str_ifneq = 'ifneq'
const token_str_ifdef = 'ifdef'
const token_str_ifndef = 'ifndef'
const token_str_else = 'else'
const token_str_endif = 'endif'
const token_str_include = 'include'
const token_str_minclude = '-include'
const token_str_colon_equals = ':='
const token_str_plus_equals = '+='
const token_str_question_equals = '?='
const token_str_equals = '='
